library verilog;
use verilog.vl_types.all;
entity AES_TOP_vlg_vec_tst is
end AES_TOP_vlg_vec_tst;
